<?xml version='1.0' encoding='UTF-8'?>

<reference anchor='I-D.ietf-anima-asa-guidelines'>
<front>
<title>Guidelines for Autonomic Service Agents</title>

<author initials='B' surname='Carpenter' fullname='Brian Carpenter'>
    <organization />
</author>

<author initials='L' surname='Ciavaglia' fullname='Laurent Ciavaglia'>
    <organization />
</author>

<author initials='S' surname='Jiang' fullname='Sheng Jiang'>
    <organization />
</author>

<author initials='P' surname='Pierre' fullname='Peloso Pierre'>
    <organization />
</author>

<date month='November' day='14' year='2020' />

<abstract><t>This document proposes guidelines for the design of Autonomic Service Agents for autonomic networks, as a contribution to describing an autonomic ecosystem.  It is based on the Autonomic Network Infrastructure outlined in the ANIMA reference model, using the Autonomic Control Plane and the Generic Autonomic Signaling Protocol.</t></abstract>

</front>

<seriesInfo name='Internet-Draft' value='draft-ietf-anima-asa-guidelines-00' />
<format type='TXT'
        target='http://www.ietf.org/internet-drafts/draft-ietf-anima-asa-guidelines-00.txt' />
</reference>
